`timescale 1ns / 1ps
//****************************************VSCODE PLUG-IN**********************************//
//----------------------------------------------------------------------------------------
// IDE :                   VSCODE     
// VSCODE plug-in version: Verilog-Hdl-Format-3.5.20250220
// VSCODE plug-in author : Jiang Percy
//----------------------------------------------------------------------------------------
//****************************************Copyright (c)***********************************//
// Copyright(C)            Please Write Company name
// All rights reserved     
// File name:              
// Last modified Date:     2025/03/11 22:50:48
// Last Version:           V1.0
// Descriptions:           
//----------------------------------------------------------------------------------------
// Created by:             Sform Chan 
// Created date:           2025/03/11 22:50:48
// mail      :             Please Write mail 
// Version:                V1.0
// TEXT NAME:              
// PATH:                   tpc
// Descriptions:           
//                         
//----------------------------------------------------------------------------------------
//****************************************************************************************//

module ysyx_25020047_IDU(
    input clk,
    input rst,
    input reg_wen,
    input  [31:0]      wdata,
    input  [31:0]       dnpc,
    input  [31:0]       inst,
    output reg [31:0]       imm,
    output reg [31:0]   inst_type,
    output [31:0]     rdata1,
    output [31:0]     rdata2,
    output [31:0]         pc,
    output [31:0]       snpc,
    output [31:0]  gpr0,
    output [31:0]  gpr1,
    output [31:0]  gpr2
);



// break down instruction

wire [6:0] opcode;
assign opcode = inst[6:0];

// Itype    
wire [4:0] Irs1;
wire [4:0] Ird;
wire [11:0] Iimm;
assign Iimm = inst[31:20];
assign Irs1 = inst[19:15];
assign Ird = inst[11:7];
wire [31:0] sIimm;
assign sIimm = {{20{Iimm[11]}}, Iimm}; // sign-extend the immediate value

// Rtype
wire [4:0] Rrs1;
wire [4:0] Rrs2;
wire [4:0] Rrd;
assign Rrd = inst[11:7];
assign Rrs1 = inst[19:15];
assign Rrs2 = inst[24:20];

// Utype
wire [4:0] Urd;
wire [19:0] Uimm;
assign Urd = inst[11:7];
assign Uimm = inst[31:12];
wire [31:0] zUimm;
assign zUimm = {Uimm, 12'b0}; // zero-extend the immediate value

// Stype
wire [4:0] Srs1;
wire [4:0] Srs2;
wire [11:0] Simm;
assign Srs1 = inst[19:15];
assign Srs2 = inst[24:20];
assign Simm = {inst[31:25], inst[11:7]};
wire [31:0] sSimm;
assign sSimm = {{20{Simm[11]}}, Simm};

// Jtype
wire [4:0] Jrd;
wire [20:0] Jimm;
assign Jimm = {inst[31], inst[19:12], inst[20], inst[30:21], 1'b0};
wire [31:0] sJimm;
assign sJimm = {{11{Jimm[20]}}, Jimm};

// Btype
wire [4:0] Brs1;
wire [4:0] Brs2;
wire [12:0] Bimm;
assign Brs1 = inst[19:15];
assign Brs2 = inst[24:20];
assign Bimm = {inst[31], inst[7], inst[30:25], inst[11:8], 1'b0};
wire [31:0] sBimm;
assign sBimm = {{19{Bimm[12]}}, Bimm};

// combine the signals
wire [4:0] rs1;
wire [4:0] rs2;
wire [4:0] rd;
assign rs1 = Rrs1 | Irs1 | Srs1 | Brs1;
assign rs2 = Rrs2 | Srs2 | Brs2;
assign rd = Rrd | Ird | Urd | Jrd;


// add more instruction types as needed  //judge the type of instruction
    always @(*)           
        begin
            casez(inst)
			//U-type
				32'b?????????????????????????0110111: inst_type = 32'h10;  // lui
				32'b?????????????????????????0010111: inst_type = 32'h200; // auipc

			//J-type
				32'b?????????????????????????1101111: inst_type = 32'h400; // jal

			//I-type	
                32'b?????????????????000?????0010011: inst_type = 32'h1; // addi
                32'b?????????????????000?????1100111: inst_type = 32'h2; // jalr
				32'b?????????????????010?????0000011: inst_type = 32'h20; // lw
                32'b?????????????????100?????0000011: inst_type = 32'h40; // lbu
				32'b?????????????????010?????0010011: inst_type = 32'h1000; //slti
				32'b?????????????????011?????0010011: inst_type = 32'h2000; //sltiu
				
			//B-type
				32'b?????????????????000?????1100011: inst_type = 32'h4000; //beq
				32'b?????????????????001?????1100011: inst_type = 32'h8000; //bne


			//R-type
                32'b00000000000100000000000001110011: inst_type = 32'h4; // ebreak
                32'b0000000??????????000?????0110011: inst_type = 32'h8; // add
				32'b0100000??????????000?????0110011: inst_type = 32'h800; // sub
				32'b0000000??????????010?????0110011: inst_type = 32'h10000; // slt
				32'b0000000??????????011?????0110011: inst_type = 32'h20000; // sltu

                
			//S-type
                32'b?????????????????010?????0100011: inst_type = 32'h80; // sw
                32'b?????????????????000?????0100011: inst_type = 32'h100; // sb
                default:                              inst_type = 32'hFFFFFFFF; // default case
            endcase                                     
        end                                          

// judge the imm
        always @(*)           
            begin                                        
                case(inst_type)
                    32'h1: imm = sIimm; // addi
                    32'h2: imm = sIimm; // jalr
					32'h20: imm = sIimm; // lw
                    32'h40: imm = sIimm; // lbu
					32'h1000: imm = sIimm; // slti
					32'h2000: imm = sIimm; // sltiu

                    32'h10: imm = zUimm; // lui
					32'h200: imm = zUimm; // auipc

                    32'h80: imm = sSimm; // sw
                    32'h100: imm = sSimm; // sb

					32'h4000: imm = sBimm; // beq
					32'h8000: imm = sBimm; // bne

					32'h400: imm = sJimm; // jal

                    default:      imm = 32'b0; // default case
                endcase
            end                                          


GPR #(5, 32) u1
(
    .clk(clk),
    .rst(rst),
    .wen(reg_wen),
    .raddr1(rs1),
    .raddr2(rs2),
    .wdata(wdata),
    .waddr(rd),
    .rdata1(rdata1),
    .rdata2(rdata2),
    .gpr0(gpr0),
    .gpr1(gpr1),
    .gpr2(gpr2)
);
 

ysyx_25020047_PC u2
(
    .clk(clk),
    .rst(rst),
    .dnpc(dnpc),
    .pc(pc),
    .snpc(snpc)
);

endmodule

